module control(instruc);

    // input     [15:0] ALU_out;
    // input     [15:0] mem_out;
    // input            mem_to_reg;

    // output    [15:0] w_data;


endmodule
module IF_ID_split();

    input            clk;
    input            rst;
    input            en;

    // data for the decode 
endmodule